module Debounce(
    input clk
     //output reg output 
);

reg previous_state;
reg [21:0]Count; //assume count is null on FPGA configuration
//--------------------------------------------
always @(posedge clk) begin
    // implement your logic here
    // button for minutes, hours and reset	 
	   // code
end 


endmodule

